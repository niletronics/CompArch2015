// =======================================================================
//   Department of Electrical and Computer Engineering
//   Portland State University
//
//   Course name:  ECE 586 - Computer Architecture
//   Term & Year:  Winter 2015
//   Instructor :  Mark Faust
//
//   Project:      PDP8 Instruction Set Architecture Simulator
//
//   Filename:     pdp.sv
// =======================================================================

`include "defines.v"
module pdp();

integer file,fileout,branchTraceFile,singleStepFile;
integer i,clk,temp1,temp2;
integer c_and,c_tad,c_isz,c_dca,c_jms,c_jmp,c_io,c_micro,c_total;	// To store counts

reg [0:31] a;
reg [0:11] PC,MQ,MB,CPMA,SR;
reg [0:11] AC;
reg [0:2]  IR;
reg        LinkBit,go,pc_inc;
reg [0:11] my_memory [0:4096];
reg [0:4]  page;
reg [0:6]  offset;
reg [0:1]  i_m;								// to store i and m bits of instruction
string     instType = "";
string     outcome = "";
reg [0:11] targetPC;
integer    int_single_step,step;
reg        step_flag = 1'b0;

//************************************************************************************** 
//********************** Register Declaration for InputOutputInst ********************** 
//**************************************************************************************
reg KCF  = 1'b0;	
reg KSF  = 1'b0;
reg KCC  = 1'b0;
reg KRS  = 1'b0;
reg KRB  = 1'b0;
reg TFL  = 1'b0;
reg TSF  = 1'b0;
reg TCF  = 1'b0;
reg TPC  = 1'b0;
reg TLS  = 1'b0;
reg SKON = 1'b0;
reg ION  = 1'b0;
reg IOF  = 1'b0;
reg KF 	 = 1'b0;
reg TF	 = 1'b0;
reg [0:7] keybuf  = 8'd0;
reg [0:7] telebuf = 8'd0; 

//************************************************************************************** 
//********************** Group 1 Microinstructions (Bit 3 = 0) ************************* 
//**************************************************************************************
reg NOP = 1'b0;					// No Operation
reg CLA = 1'b0;					// CLear Accumulator (1)
reg CLL = 1'b0;					// CLear Link (1)
reg CMA = 1'b0;					// Complement Accumulator (2)
reg CML = 1'b0;					// Complement Link (2)
reg IAC = 1'b0;					// Increment ACumulator (3)
reg RAR = 1'b0;					// Rotate Accumulator and link Right (4)
reg RTR = 1'b0;					// Rotate accumulator and link Right Twice (4)
reg RAL = 1'b0;					// Rotate Accumulator and link Left (4)
reg RTL = 1'b0;					// Rotate Accumulator and link left Twice (4)

//************************************************************************************** 
//*************** Group 2 Microinstructions (Bit 3 = 1, Bit 11 = 0) ********************
//**************************************************************************************
reg SMA = 1'b0;					// Skip on Minus Accumulator (1)
reg SZA = 1'b0;					// Skip on Zero Accumulator (1)
reg SNL = 1'b0;					// Skip on Nonzero Link (1)
reg SPA = 1'b0;					// Skip on Positive Accumulator (1)
reg SNA = 1'b0;					// Skip on Nonzero Accumulator (1)
reg SZL = 1'b0;					// Skip on Zero Link (1)
reg SKP = 1'b0;					// SkiP always (1)
reg OSR = 1'b0;					// Or Switch Register with accumulator (3)
reg HLT = 1'b0;					// Halt (3)

//************************************************************************************** 
//*************** Group 3 Microinstructions (Bit 3 = 1, Bit 11 = 1) ********************
//**************************************************************************************
reg MQL = 1'b0;					// Load MQ register from AC and Clear AC (2); C(MQ) <- C(AC); C(AC) <- 0;
reg MQA = 1'b0;					// Or AC with MQ register (2) ; C(AC) <- C(AC) Or C(MQ)
reg SWP = 1'b0;					// Swap AC and MQ registers (3)
reg CAM = 1'b0;					// Clear AC and MQ registers (3)
reg ORSubgroup  = 1'b0;				// Condition for ORSubGroup 1'b1 = True, 1'b0 = False
reg ANDSubgroup = 1'b0;				// Condition for ANDSubgroup  1'b1 = True, 1'b0 = False

reg int_JMS = 1'b0;				// JMS flag for Branch Trace File
reg int_JMP = 1'b0;				// JMP flag for Branch Trace File
reg int_ISZ = 1'b0;				// ISZ flag for Branch Trace File
reg [0:15] single_step;

parameter AND = 3'd0,				// Memory reference instructions
	  TAD = 3'd1,
	  ISZ = 3'd2, 
	  DCA = 3'd3,
	  JMS = 3'd4,
	  JMP = 3'd5,
	  IO  = 3'd6,
	  M_INSTRUCTIONS = 3'd7,

	  i_KCF = 12'o6030,			// Clear Keyboard Flag
      	  i_KSF = 12'o6031,			// Skip on Keyboard Flag set
      	  i_KCC = 12'o6032,			// Clear Keyboard flag and ACC
      	  i_KRS = 12'o6034,			// Read Keyboard buffer Static A
      	  i_KRB = 12'o6036,			// Read Keyboard Buffer dynamic 

//*********************** Printer (CRT) - Device #4 **************************
      	  i_TFL = 12'o6040,			// Set printer flag
     	  i_TSF = 12'o6041,			// Skip on printer flag set
      	  i_TCF = 12'o6042,			// Clear printer Flag
      	  i_TPC = 12'o6044,			// Load printer buffer with ACC
      	  i_TLS = 12'o6046,			// Load printer Sequence ; Print

//*********************** Interrupt System - Device #0 ***********************
       	  i_SKON = 12'o6000,			// Skip if the interrupt system 
      	  i_ION  = 12'o6001,			// Execute the next instruction 
      	  i_IOF  = 12'o6002,			// Turn the interrupt system off

//**************************** Group 3 instructions ***************************
	  i_CLA = 12'o7601,
	  i_MQL = 12'o7421, 
	  i_MQA = 12'o7501,
	  i_SWP = 12'o7521,
	  i_CAM = 12'o7621;

//=============================================================================
//=============================================================================

initial 
begin
$display("********************* ISA SIMULATOR *********************");
initializeVariables();
initialize();
page=PC[0:4];
offset=PC[5:11];
go=1'b1;

	fileout=$fopen("output.txt","w");
	branchTraceFile=$fopen("Branch_Trace.txt","w");
	$fwrite(branchTraceFile,"CURRENT PC \t INSTRUCTION \t TARGET PC \t BRANCH OUTCOME \n");
	$fwrite(branchTraceFile,"---------------------------------------------------------------\n");
	$display("Do you want single stepping? Y/N (y/n) :");
	step = $fgetc('h8000_0000);

	while(go==1'b1&&PC!=`EOMemory)
	begin
		if(step == "Y" || step == "y")
		begin
			$display("Press any key to continue \n");		// Single stepping. Press ENTER to continue
			int_single_step = $fgetc('h8000_0000);
			step_flag = 1'b1;
			
		end

		pc_inc=0;
		MemoryRead(`instruction);// 0 indicates that we are fetching instruction and we write 1 when we want data
		int_JMS = 1'b0;
		int_JMP = 1'b0;
		int_ISZ = 1'b0;
		SMA = 1'b0;					
		SZA = 1'b0;				
		SNL = 1'b0;					
		SPA = 1'b0;					
		SNA = 1'b0;					
		SZL = 1'b0;					
		SKP = 1'b0;	
		KSF = 1'b0;
		TSF = 1'b0;	

		case(IR)
	   	AND: begin
			c_and=c_and+1;
			effectiveAddress();	// to calculate effective address
			MemoryRead(`data);	// to get the contents of effective address
			AC=AC&MB;
			clk=clk+2;
			//`ifdef SHOW
			//$display("PC is %o and AC is %o",PC,AC);
			//`endif
			if(step_flag) begin $display("AND"); end
		     end

	   	TAD: begin
			c_tad=c_tad+1;
			effectiveAddress();	// to calculate effective address
			MemoryRead(`data);
			if((AC < 12'd2048 && MB < 12'd2048 &&(AC+MB) > 12'd2047)||(AC > 12'd2047 && MB > 12'd2047 &&(AC+MB) < 12'd2048))
		    		$display("Overflow occured");
			{LinkBit,AC}={LinkBit,AC}+MB;
			clk=clk+2;
			//`ifdef SHOW
			//$display("PC is %o and AC is %o",PC,AC);
			//`endif
			if(step_flag) begin $display("TAD"); end
		     end

	   	ISZ: begin
			c_isz=c_isz+1;
			effectiveAddress();	// to calculate effective address
			MemoryRead(`data);
			MB=MB+1;
			MemoryWrite(MB);
			if(MB==0)
		    		pc_inc=1'b1;			//FLAG FOR PC=PC+1;
			clk=clk+2;
			int_ISZ = 1'b1;
			if(step_flag) begin $display("ISZ"); end
		     end

	   	DCA: begin
			c_dca=c_dca+1;
			effectiveAddress();	// to calculate effective address
			MemoryWrite(AC);
			AC=0;
			clk=clk+2;
			if(step_flag) begin $display("DCA"); end
		     end
	   	JMS: begin
	   		c_jms=c_jms+1;
			effectiveAddress();	
			MemoryWrite(PC+1);
			clk=clk+2;
			int_JMS = 1'b1;
			if(step_flag) begin $display("JMS"); end
		     end

	   	JMP: begin
			c_jmp=c_jmp+1;
			effectiveAddress();		
			clk=clk+1;
			int_JMP = 1'b1;
			if(step_flag) begin $display("JMP"); end
		     end

	   	IO: begin
			c_io=c_io+1;
			InputOutputInst();
			if(step_flag) begin $display("IO"); end
		    end

	   	M_INSTRUCTIONS: begin
			c_micro=c_micro+1;
			if(i_m[0]==0)
		   		Group1MicroInstructions();
			else if(i_m[0]==1&&offset[6]==0)
		   		Group2MicroInstructions();
			else if(i_m[0]==1&&offset[6]==1)
		   		Grp3MicroInstruction();
			clk=clk+1;
		    end
		endcase

		if(step_flag)
		begin
			$display("In octal PC: %o \t AC: %o \t LinkBit: %o ",PC,AC,LinkBit);
		end
		branchTrace();

		if(IR==JMS) 	 begin PC=CPMA+1; end		// Write return address
		else if(IR==JMP) begin PC=CPMA;   end			
		else if(pc_inc==1'b1)	begin PC=PC+2;   end
		else PC=PC+1;
	end


$display("\n***************************************************"); 
$display("********************* SUMMARY *********************"); 
$display("***************************************************\n"); 
summary();

$fclose(fileout);
$fclose(branchTraceFile);
end

//========================================================================================================
//========================================= Summary ======================================================
//========================================================================================================
task summary;
begin
c_total= c_and+c_tad+c_isz+c_dca+c_jms+c_jmp+c_io+c_micro;
$display("No. of AND instructions :    \t %d",c_and);
$display("No. of TAD instructions :    \t %d",c_tad);
$display("No. of ISZ instructions :    \t %d",c_isz);
$display("No. of DCA instructions :    \t %d",c_dca);
$display("No. of JMS instructions :    \t %d",c_jms);
$display("No. of JMP instructions :    \t %d",c_jmp);
$display("No. of IO instructions :     \t %d",c_io);
$display("No. of MICRO instructions :  \t %d",c_micro);
$display("No. of TOTAL instructions :  \t %d",c_total);
$display("Total clock cycles required :\t %d",clk);
$display("PC IS %o",PC);
$display("Accumulator:%o and LinkBit:%o",AC,LinkBit);
end

endtask

//========================================================================================================
//========================================= Variable initialization ======================================
//========================================================================================================
task initializeVariables;
begin
a=0;
clk=0;
c_and=0;c_tad=0;c_isz=0;c_dca=0;c_jms=0;c_jmp=0;c_io=0;c_micro=0;c_total=0;pc_inc=0;
step_flag=1'b0;
AC=12'b0;
LinkBit=1'b0;
end
endtask
//========================================================================================================
//========================================= Address Calculation ==========================================
//========================================================================================================
task intaddress;
input [0:31]a1;
output decaddr;
integer decaddr,x,y,z,flag,address;
begin
	flag=0;
	if(a1[8:15]>47&&a1[8:15]<58)
		x=48;
	else if(a1[8:15]>64&&a1[8:15]<71)
		x=55;
	else if(a1[8:15]>96&&a1[8:15]<103)
		x=87;
	else
		flag=1;
	if(a1[16:23]>47&&a1[16:23]<58)
		y=48;
	else if(a1[16:23]>64&&a1[16:23]<71)
		y=55;
	else if(a1[16:23]>96&&a1[16:23]<103)
		y=87;
	else
		flag=1;
	if(a1[24:31]>47&&a1[24:31]<58)
		z=48;
	else if(a1[24:31]>64&&a1[24:31]<71)
		z=55;
	else if(a1[24:31]>96&&a1[24:31]<103)
		z=87;
	else
		flag=1;

if(flag==0)
	begin
	decaddr=((a1[8:15]-x)*256)+((a1[16:23]-y)*16)+(a1[24:31]-z);
	//$display("dec address %d",decaddr);
	end
else
	decaddr=5000;// not a vaild address.
	
end
endtask

//========================================================================================================
//============================================= Initialize ===============================================
//========================================================================================================

task initialize;
integer temp,b;
reg [500*8-1:0] file_name;
begin
$display("Enter file name :");
b = $fgets(file_name, 'h8000_0000);
file_name = file_name >> 8;

file = $fopen(file_name,"r");
// checking if file is not empty or invalid
if(file == `NULL) 
	begin
	$display("Error reading file");
	end
else 
	begin	
	$readmemh(file_name, my_memory);
	/*for(i=0;i<4095;i=i+1)  // to display contents of memory
	   begin
	   if(my_memory[i]!==12'hxxx)
           $display("%d %h",i,my_memory[i]);
	   end*/
	b=$fscanf(file,"%s",a);
	if(a[0:7]=="@")
	   begin
	   $display("yes");
	   intaddress(a,temp);
	   if(temp!=5000)
	      PC=temp;
	   else
	      $display("Invalid Address");
	   end
	else
	   PC=128;
	end
$display("PC is %d",PC);
$fclose(file_name);

// initialize keyboard buffer with random value and set KF flag
// mimic the keyboard input :-)
keybuf	= $random;
//keybuf = 8'd7;
KF	= 1'b1;
TF = 1'b1;
end
endtask

//========================================================================================================
//=================================== EffectiveAddress Calculation =======================================
//========================================================================================================

task effectiveAddress;
begin
if(i_m==2'b00)
	CPMA={5'b00000,offset};
else if(i_m==2'b01)
	CPMA={page,offset};
else if(i_m[0]==1)
	begin
	clk=clk+1;
	if(offset>7'b0000111 && offset < 7'b0010000 && i_m[1]==0)
	   begin
		    clk=clk+1;
	            CPMA= my_memory[{5'b00000,offset}]+1; // removed 1 my_memory 
		    my_memory[{5'b00000,offset}]=my_memory[{5'b00000,offset}]+1;// confirm correctness.
		    $fwrite(fileout,"%d %o \n",0,{5'b00000,offset});
		    $fwrite(fileout,"%d %o \n",1,{5'b00000,offset});		    
		 
           end
        else
	   begin
		if(i_m[1]==0)
		    begin
		    CPMA=my_memory[{5'b00000,offset}];// 2 memory references for these 
	            $fwrite(fileout,"%d %o \n",0,{5'b00000,offset});
                    end
		else
		    begin
		    CPMA=my_memory[{page,offset}];// 2 memory references for these 
	            $fwrite(fileout,"%d %o \n",0,{page ,offset});
		    end
	   end
	end
end
endtask

//========================================================================================================
//============================================ Memory Read ===============================================
//========================================================================================================

task MemoryRead;
input i;
integer i;

begin
	if(i==0)				// Instruction fetch
	begin
        	IR=my_memory[PC][0:2];
		i_m=my_memory[PC][3:4];
		offset=my_memory[PC][5:11];	// This offset will be used in effective address calculation
		page=PC[0:4];
	 	$fwrite(fileout,"%d %o \n",2,PC);
	end
	else
	begin
		MB=my_memory[CPMA];
		$fwrite(fileout,"%d %o \n",0,CPMA);
	end
end
endtask

//========================================================================================================
//============================================ Memory Write ==============================================
//========================================================================================================

task MemoryWrite;
input reg [0:11] out_data; 
begin
	MB=out_data;
	my_memory[CPMA]=MB;
	$fwrite(fileout,"%d %o \n",1,CPMA);
end
endtask

//========================================================================================================
//====================================== Input Output Instructions =======================================
//========================================================================================================

task InputOutputInst;

integer IO_char_handler;
reg [500*8-1:0] IO_char;

begin

if(my_memory[PC] == i_KCF) begin KCF =1'b1; if(step_flag) begin $display("KCF "); end end else KCF = 1'b0;
if(my_memory[PC] == i_KSF) begin KSF =1'b1; if(step_flag) begin $display("KSF "); end end else KSF = 1'b0;
if(my_memory[PC] == i_KCC) begin KCC =1'b1; if(step_flag) begin $display("KCC "); end end else KCC = 1'b0;
if(my_memory[PC] == i_KRS) begin KRS =1'b1; if(step_flag) begin $display("KRS "); end end else KRS = 1'b0;
if(my_memory[PC] == i_KRB) begin KRB =1'b1; if(step_flag) begin $display("KRB "); end end else KRB = 1'b0;
                         
if(my_memory[PC] == i_TFL) begin TFL =1'b1; if(step_flag) begin $display("TFL "); end end else TFL = 1'b0;
if(my_memory[PC] == i_TSF) begin TSF =1'b1; if(step_flag) begin $display("TSF "); end end else TSF = 1'b0;
if(my_memory[PC] == i_TCF) begin TCF =1'b1; if(step_flag) begin $display("TCF "); end end else TCF = 1'b0;
if(my_memory[PC] == i_TPC) begin TPC =1'b1; if(step_flag) begin $display("TPC "); end end else TPC = 1'b0;
if(my_memory[PC] == i_TLS) begin TLS =1'b1; if(step_flag) begin $display("TLS "); end end else TLS = 1'b0;
                         
if(my_memory[PC]== i_SKON) begin SKON=1'b1; if(step_flag) begin $display("SKON"); end end else SKON = 1'b0;
if(my_memory[PC] == i_ION) begin ION =1'b1; if(step_flag) begin $display("ION "); end end else ION = 1'b0;
if(my_memory[PC] == i_IOF) begin IOF =1'b1; if(step_flag) begin $display("IOF "); end end else IOF = 1'b0;

	// INPUT

	if(KCF) KF = 1'b0;
	if(KSF && KF) begin pc_inc = 1'b1; end

	if(KCC) 
	begin
		KF = 1'b0;
		AC = 12'b0;
	end

	if(KRS)
	begin
		$display("Enter a character from keyboard :");
		$fflush('h8000_0000);
		IO_char_handler = $fgetc('h8000_0000);
		if(!step_flag) begin IO_char_handler = $fgetc('h8000_0000); end
		keybuf = IO_char_handler;
		if(step_flag) begin $display("KRS : %c", keybuf); end
		AC[4:11] |= keybuf;
	end

	if(KRB)
	begin
		$display("Enter a character from keyboard :");
		$fflush('h8000_0000);
		IO_char_handler = $fgetc('h8000_0000);
		if(!step_flag) begin IO_char_handler = $fgetc('h8000_0000); end
		keybuf = IO_char_handler;
		if(step_flag) begin $display("KRB : %c", keybuf); end
		AC = {4'h0,keybuf};
		KF = 1'b0;
	end

	//OUTPUT

	if(TFL) TF = 1'b1;
	if(TSF && TF) pc_inc = 1'b1; 
	if(TCF) TF = 1'b0;

	if(TPC) 
	begin
		telebuf = AC[4:11];
		$display("*********************");
		$display("PRINTER OUTPUT => \"%c\"",telebuf);
		$display("*********************");
	end

	if(TLS)
	begin
		telebuf = AC[4:11];
		TF = 1'b0;
		$display("*********************");
		$display("PRINTER OUTPUT => \"%c\"",telebuf);
		$display("*********************");
	end                                   
end
endtask

//========================================================================================================
//======================================= Group 2 Microinstructions ======================================
//========================================================================================================

task Group2MicroInstructions;  
static integer Grp2Cnt;
begin
//	if(my_memory[PC] ==? 12'b111_1?0_001_??0) begin	SKP	=1'b1; $display("SKP"); end else SKP	=1'b0;
//	if(my_memory[PC] ==? 12'b111_11?_???_??0) begin	CLA	=1'b1; $display("CLA"); end else CLA	=1'b0;
//	if(my_memory[PC] ==? 12'b111_1??_???_1?0) begin	OSR	=1'b1; $display("OSR"); end else OSR	=1'b0;
//	if(my_memory[PC] ==? 12'b111_1??_???_?10) begin	HLT	=1'b1; $display("HLT"); end else HLT	=1'b0;
//	if(my_memory[PC] ==? 12'b111_1?1_??0_??0) begin	SMA	=1'b1; $display("SMA"); end else SMA	=1'b0;
//	if(my_memory[PC] ==? 12'b111_1??_1?0_??0) begin	SZA	=1'b1; $display("SZA"); end else SZA	=1'b0;
//	if(my_memory[PC] ==? 12'b111_1??_?10_??0) begin	SNL	=1'b1; $display("SNL"); end else SNL	=1'b0;
//	if(my_memory[PC] ==  12'b111_100_000_000) begin	NOP	=1'b1; $display("NOP"); end else NOP	=1'b0;
//	if(my_memory[PC] ==? 12'b111_1?1_??1_??0) begin	SPA	=1'b1; $display("SPA"); end else SPA	=1'b0;
//	if(my_memory[PC] ==? 12'b111_1??_1?1_??0) begin	SNA	=1'b1; $display("SNA"); end else SNA	=1'b0;
//	if(my_memory[PC] ==? 12'b111_1??_?11_??0) begin	SZL	=1'b1; $display("SZL"); end else SZL	=1'b0;

	if(my_memory[PC] ==? 12'b111_1?0_001_??0) begin	SKP	=1'b1; if(step_flag) begin $display("SKP"); end end else SKP	=1'b0;
	if(my_memory[PC] ==? 12'b111_11?_???_??0) begin	CLA	=1'b1; if(step_flag) begin $display("CLA"); end end else CLA	=1'b0;
	if(my_memory[PC] ==? 12'b111_1??_???_1?0) begin	OSR	=1'b1; if(step_flag) begin $display("OSR"); end end else OSR	=1'b0;
	if(my_memory[PC] ==? 12'b111_1??_???_?10) begin	HLT	=1'b1; if(step_flag) begin $display("HLT"); end end else HLT	=1'b0;
	if(my_memory[PC] ==? 12'b111_1?1_??0_??0) begin	SMA	=1'b1; if(step_flag) begin $display("SMA"); end end else SMA	=1'b0;
	if(my_memory[PC] ==? 12'b111_1??_1?0_??0) begin	SZA	=1'b1; if(step_flag) begin $display("SZA"); end end else SZA	=1'b0;
	if(my_memory[PC] ==? 12'b111_1??_?10_??0) begin	SNL	=1'b1; if(step_flag) begin $display("SNL"); end end else SNL	=1'b0;
	if(my_memory[PC] ==  12'b111_100_000_000) begin	NOP	=1'b1; if(step_flag) begin $display("NOP"); end end else NOP	=1'b0;
	if(my_memory[PC] ==? 12'b111_1?1_??1_??0) begin	SPA	=1'b1; if(step_flag) begin $display("SPA"); end end else SPA	=1'b0;
	if(my_memory[PC] ==? 12'b111_1??_1?1_??0) begin	SNA	=1'b1; if(step_flag) begin $display("SNA"); end end else SNA	=1'b0;
	if(my_memory[PC] ==? 12'b111_1??_?11_??0) begin	SZL	=1'b1; if(step_flag) begin $display("SZL"); end end else SZL	=1'b0;
	//Condition checking for SubGroup
	if((SMA && AC[0]==1'b1) || (SZA && AC == 12'b0) || (SNL && LinkBit==1'b1)) ORSubgroup =1'b1; else ORSubgroup =1'b0;
	
	if(SPA || SNA || SZL )	begin
		if(((SPA && AC[0]==1'b0) || !SPA) && ((SNA && AC != 12'b0)||!SNA) && ((SZL && LinkBit==1'b0)||!SZL)) 
			ANDSubgroup =1'b1; 
		else 
			ANDSubgroup =1'b0;
	end
	else
	ANDSubgroup =1'b0;	
	
	if(ORSubgroup || ANDSubgroup || SKP) pc_inc = 1'b1; 					//OR SubGroup, later combining common case						// Priority(1)
	if(CLA) AC = 12'b0;						// Priority (2)
	if(OSR) AC = (AC | SR);						// Priority (3)
	if(NOP) $display("NOP is encounter at PC = %h and Memory= %o",PC,my_memory[PC]);
	if(HLT) go = 1'b0;						// Priority (3) //Assuming HLT should be executed as the last instruction 
	
	if(SKP||CLA||OSR||HLT||SMA||SZA||SNL||NOP||SPA||SNA||SZL)
		Grp2Cnt++;
	else 
		$display("Invalid Group2MicroInstructions : Instruction = %o and PC = %d",my_memory[PC],PC);
end
endtask

//========================================================================================================
//======================================= Group 1 Microinstructions ======================================
//========================================================================================================

task Group1MicroInstructions;
reg LinkBitLocal;
begin
if(my_memory[PC] ==? 12'b111_000_000_000) begin NOP = 1'b1;	if(step_flag) $display("NOP"); end else NOP =1'b0;
if(my_memory[PC] ==? 12'b111_01?_???_???) begin CLA = 1'b1;	if(step_flag) $display("CLA"); end else CLA =1'b0;
if(my_memory[PC] ==? 12'b111_0?1_???_???) begin CLL = 1'b1;	if(step_flag) $display("CLL"); end else CLL =1'b0;
if(my_memory[PC] ==? 12'b111_0??_1??_???) begin CMA = 1'b1;	if(step_flag) $display("CMA"); end else CMA =1'b0;
if(my_memory[PC] ==? 12'b111_0??_?1?_???) begin CML = 1'b1;	if(step_flag) $display("CML"); end else CML =1'b0;
if(my_memory[PC] ==? 12'b111_0??_???_??1) begin IAC = 1'b1;	if(step_flag) $display("IAC"); end else IAC =1'b0;
if(my_memory[PC] ==? 12'b111_0??_??1_?0?) begin RAR = 1'b1;	if(step_flag) $display("RAR"); end else RAR =1'b0;
if(my_memory[PC] ==? 12'b111_0??_???_10?) begin RAL = 1'b1;	if(step_flag) $display("RAL"); end else RAL =1'b0;
if(my_memory[PC] ==? 12'b111_0??_??1_?1?) begin RTR = 1'b1;	if(step_flag) $display("RTR"); end else RTR =1'b0;
if(my_memory[PC] ==? 12'b111_0??_???_11?) begin RTL = 1'b1;	if(step_flag) $display("RTL"); end else RTL =1'b0;

	if(NOP) $display("NOP ENCOUNTERED AT PC = %o and my_memory[PC]=%o",PC,my_memory[PC]);
	if(CLA) 
	begin
		AC = 12'b0;        // priority_1
 		//$display("CLA Executed CLA = %o", AC);
		if(step_flag) 
		begin 
			$display("CLA Executed CLA = %o", AC); 
		end
        end

if(CLL) LinkBit = 1'b0;

if(CMA) AC = ~AC;          // priority_2
if(CML) LinkBit = ~LinkBit;

	if(IAC) 
	begin	
    		if((AC+1)>12'd2047&&AC < 12'd2048)
    		begin
    			$display("Overflow occured");
    		end
    		{LinkBit,AC}={LinkBit,AC}+1'b1;

end

	if(RAR) 
	begin 
		if(step_flag) begin $display("RAR Executed AC Pre = %o", AC); end
		LinkBitLocal = AC [11]; 
		AC = {LinkBit,AC[0:10]};
		LinkBit = LinkBitLocal; 
		if(step_flag) begin $display("RAR Executed AC Aftervalue = %o", AC); end 
	end  //priority_4

if(RAL) begin 
	if(step_flag) begin $display("RAL Executed AC Pre = %o", AC); end
	LinkBitLocal = AC [0];  
	AC = {AC[1:11],LinkBit};
	LinkBit = LinkBitLocal; 
	if(step_flag) begin $display("CLA Executed AC Aftervalue = %o", AC); end
end
              
if(RTR) begin 
	if(step_flag) begin $display("RTR Executed AC Pre = %o", AC); end
	LinkBitLocal = AC[10];
	AC = {AC[11], LinkBit, AC[0:9]};
	LinkBit = LinkBitLocal;
end //priority_5

if(RTL) begin
	if(step_flag) begin $display("RTL Executed AC Pre = %o", AC); end
	LinkBitLocal = AC[1]; 
	AC = {AC[2:11], LinkBit, AC[0]};
	LinkBit = LinkBitLocal;
end   

end
endtask


//========================================================================================================
//======================================= Group 3 Microinstructions ======================================
//========================================================================================================

task Grp3MicroInstruction();
begin
	integer Grp3Cnt;
	if(my_memory[PC] == i_CLA ) begin	CLA =1'b1; if(step_flag) begin $display("CLA"); end end else CLA = 1'b0;
	if(my_memory[PC] == i_MQL ) begin	MQL =1'b1; if(step_flag) begin $display("MQL"); end end else MQL = 1'b0;
	if(my_memory[PC] == i_MQA ) begin	MQA =1'b1; if(step_flag) begin $display("MQA"); end end else MQA = 1'b0;
	if(my_memory[PC] == i_SWP ) begin	SWP =1'b1; if(step_flag) begin $display("SWP"); end end else SWP = 1'b0;
	if(my_memory[PC] == i_CAM ) begin	CAM =1'b1; if(step_flag) begin $display("CAM"); end end else CAM = 1'b0;

	if(CLA) AC = 12'b0;	
	if(MQL) 
	begin 
		MQ [0:11] =  AC[0:11];
		AC [0:11] = 12'b0;
	end
	if (MQA) AC = AC | MQ;
	if (SWP) 
	begin
		MQ <= AC;
		AC <= MQ;
	end
	if (CAM) 
	begin
		AC [0:11] = 12'b0;
		MQ [0:11] = 12'b0;
	end

if(CLA || MQL || MQA || SWP || CAM )
	Grp3Cnt++;
else 
	$display("Invalid Group 3 MircoInstruction at PC = %d \n Instruction = %o", PC, my_memory[PC]);
end
if(step_flag) begin
	$display("AC = %o, MQ = %o, LinkBit = %b, PC = %d ",AC,MQ,LinkBit,PC);
end 
		
endtask

//========================================================================================================
//=========================================== Branch Trace File ==========================================
//========================================================================================================

task branchTrace();
begin
	instType = "";

	case({SMA,SZA,SNL})
		3'b111 : instType = "SMA SZA SNL";
		3'b110 : instType = "SMA SZA";
		3'b101 : instType = "SMA SNL";
		3'b100 : instType = "SMA";
		3'b011 : instType = "SZA SNL";
		3'b010 : instType = "SZA";
		3'b001 : instType = "SNL";
	endcase

	case({SPA,SNA,SZL})
		3'b111 : instType = "SPA,SNA,SZL";
		3'b110 : instType = "SPA SNA";
		3'b101 : instType = "SPA SZL";
		3'b100 : instType = "SPA";
		3'b011 : instType = "SNA SZL";
		3'b010 : instType = "SNA";
		3'b001 : instType = "SZL";
	endcase

	if(SKP == 1)   begin instType = "SKP"; end
	if(int_JMP == 1) begin instType = "JMP"; end
	if(int_JMS == 1) begin instType = "JMS"; end
	if(int_ISZ == 1)   begin instType = "ISZ"; end
	if(KSF) begin instType = "KSF"; end
	if(TSF) begin instType = "TSF"; end

	if(int_JMP || int_JMS || pc_inc) begin 
		outcome = "TAKEN"; 
	end
	else begin 
		outcome = "NOT TAKEN"; 
	end

	if(pc_inc) begin 
		targetPC = PC + 2; 
	end
	else if(int_JMP) begin 
		targetPC = CPMA;
	end
	else if(int_JMS) begin 
		targetPC = CPMA + 1'b1;  
	end
	else if(SMA || SZA || SNL || SPA || SNA || SZL || ISZ || KSF || TSF) begin
		targetPC = PC + 1;
	end

	if(SMA || SZA || SNL || SPA || SNA || SZL || SKP || int_ISZ || KSF || TSF)
	begin
		$fwrite(branchTraceFile,"%8o \t %8s \t %8o \t %8s \n",PC,instType,targetPC,outcome);
	end
	else if (int_JMP || int_JMS)
	begin
		$fwrite(branchTraceFile,"%8o \t %8s \t %8o \t %8s \n",PC,instType,targetPC,outcome);
	end
end
endtask
endmodule
