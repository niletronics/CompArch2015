task MemoryRefJMP;
begin
	effectiveAddress();	
end
endtask

