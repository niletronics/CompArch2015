task MemoryRefJMS;
begin
	effectiveAddress();	
	MemoryWrite(PC+1);
end
endtask

