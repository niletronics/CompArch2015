`include "defines.v"

module pdp8(); //Signals listing for testbench




endmodule