`include "defines.v"

module pdp8_tb();

endmodule
